
interface ltssm_if(input logic clk);
    logic rst_n;
    logic valid;
    logic [31:0] ts_data;
endinterface
